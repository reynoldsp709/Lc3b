library verilog;
use verilog.vl_types.all;
entity memory_test is
end memory_test;
