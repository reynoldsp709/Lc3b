library verilog;
use verilog.vl_types.all;
entity shift_test is
end shift_test;
