library verilog;
use verilog.vl_types.all;
entity regfile_test is
end regfile_test;
