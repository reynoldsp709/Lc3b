library verilog;
use verilog.vl_types.all;
entity gate_test is
end gate_test;
