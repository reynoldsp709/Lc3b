library verilog;
use verilog.vl_types.all;
entity zext_test is
end zext_test;
